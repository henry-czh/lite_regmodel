
package lite_regmodel;
    `include "lite_reg_macros.svh"
    `include "dpi/uvm_hdl.svh"
    `include "dpi/uvm_svcmd_dpi.svh"
    `include "dpi/uvm_regex.svh"
    `include "lite_adaptor.sv"
    `include "lite_field.sv"
    `include "lite_reg.sv"
    `include "lite_regmodel.sv"
    `include "lite_reset_check_tc.sv"
    `include "lite_hdl_path_check_tc.sv"
    `include "lite_access_check_tc.sv"
endpackage

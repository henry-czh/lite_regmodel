
class lite_regmodel;
endclass


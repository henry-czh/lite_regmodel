
class lite_regmodel;
    function new(string name="");
        
    endfunction
endclass

